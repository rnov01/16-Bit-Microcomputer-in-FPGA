
module pll (
	clk_25_clk,
	clk_in_clk,
	rst_reset);	

	output		clk_25_clk;
	input		clk_in_clk;
	input		rst_reset;
endmodule
