-- pll.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pll is
	port (
		clk_25_clk : out std_logic;        -- clk_25.clk
		clk_in_clk : in  std_logic := '0'; -- clk_in.clk
		rst_reset  : in  std_logic := '0'  --    rst.reset
	);
end entity pll;

architecture rtl of pll is
	component pll_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component pll_video_pll_0;

begin

	video_pll_0 : component pll_video_pll_0
		port map (
			ref_clk_clk        => clk_in_clk, --      ref_clk.clk
			ref_reset_reset    => rst_reset,  --    ref_reset.reset
			vga_clk_clk        => clk_25_clk, --      vga_clk.clk
			reset_source_reset => open        -- reset_source.reset
		);

end architecture rtl; -- of pll
